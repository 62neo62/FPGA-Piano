//utilizing decimal representation for half period clock cycles

timescale 1 ns / 1 ps
// Declare the module and its ports. This is
// using Verilog-2001 syntax.
module piano (
 input wire clk,
 input wire hush,
 input wire [3:0] note,
 output wire speaker
 );

reg

case @*
val = 17'd113635;
        4'b0001:
        val = 17'd107257;
        4'b0010:
        val = 17'd101237;
        4'b0011:
        val = 17'd95555;
        4'b0100:
        val = 17'd90192;
        4'b0101:
        val = 17'd85130;
        4'b0110:
        val = 17'd80352;
        4'b0111:
        val = 17'd75842;
        4'b1000:
        val = 17'd71585;
        4'b1001:
        val = 17'd67568;
        4'b1010:
        val = 17'd63775;
        4'b1011:
        val = 17'd60196;
        4'b1100:
        val = 17'd56817;
        4'b1101:
        val = 17'd53628;
        4'b1110:
        val = 17'd50618;
        4'b1111:
        val = 17'd47777;
endmodule

initial
begin
	speakeractive <= 0;
	counter <=0:
end
always(posedge clk)
begin
	counter <=0;
	speakeractive <= outclock;
	if((counter == frequency) && (hush == 1'b0)) //counter is equal to freq and hush/mute not pressed
	begin
		counter <=0;
		speakeractive <= !speakeractive;
	end
end
	endmodule
